// nios2_qsys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios2_qsys (
		input  wire        clk_clk,       //     clk.clk
		output wire        epcs_dclk,     //    epcs.dclk
		output wire        epcs_sce,      //        .sce
		output wire        epcs_sdo,      //        .sdo
		input  wire        epcs_data0,    //        .data0
		input  wire [3:0]  key_export,    //     key.export
		output wire [3:0]  led_export,    //     led.export
		input  wire        reset_reset_n, //   reset.reset_n
		output wire [10:0] sdram47_addr,  // sdram47.addr
		output wire [1:0]  sdram47_ba,    //        .ba
		output wire        sdram47_cas_n, //        .cas_n
		output wire        sdram47_cke,   //        .cke
		output wire        sdram47_cs_n,  //        .cs_n
		inout  wire [31:0] sdram47_dq,    //        .dq
		output wire [3:0]  sdram47_dqm,   //        .dqm
		output wire        sdram47_ras_n, //        .ras_n
		output wire        sdram47_we_n   //        .we_n
	);

	wire  [31:0] nios2_data_master_readdata;                                  // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                               // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                               // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [23:0] nios2_data_master_address;                                   // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                                      // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_readdatavalid;                             // mm_interconnect_0:nios2_data_master_readdatavalid -> nios2:d_readdatavalid
	wire         nios2_data_master_write;                                     // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                 // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                           // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [23:0] nios2_instruction_master_address;                            // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                               // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire         nios2_instruction_master_readdatavalid;                      // mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;            // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;         // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;         // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;             // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;          // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;               // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;           // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_epcs_control_port_chipselect;         // mm_interconnect_0:epcs_epcs_control_port_chipselect -> epcs:chipselect
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_readdata;           // epcs:readdata -> mm_interconnect_0:epcs_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_epcs_control_port_address;            // mm_interconnect_0:epcs_epcs_control_port_address -> epcs:address
	wire         mm_interconnect_0_epcs_epcs_control_port_read;               // mm_interconnect_0:epcs_epcs_control_port_read -> epcs:read_n
	wire         mm_interconnect_0_epcs_epcs_control_port_write;              // mm_interconnect_0:epcs_epcs_control_port_write -> epcs:write_n
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_writedata;          // mm_interconnect_0:epcs_epcs_control_port_writedata -> epcs:writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                         // mm_interconnect_0:ram_s1_chipselect -> ram:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                           // ram:readdata -> mm_interconnect_0:ram_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                            // mm_interconnect_0:ram_s1_address -> ram:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                         // mm_interconnect_0:ram_s1_byteenable -> ram:byteenable
	wire         mm_interconnect_0_ram_s1_write;                              // mm_interconnect_0:ram_s1_write -> ram:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                          // mm_interconnect_0:ram_s1_writedata -> ram:writedata
	wire         mm_interconnect_0_ram_s1_clken;                              // mm_interconnect_0:ram_s1_clken -> ram:clken
	wire  [31:0] mm_interconnect_0_pio_key_s1_readdata;                       // pio_key:readdata -> mm_interconnect_0:pio_key_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_key_s1_address;                        // mm_interconnect_0:pio_key_s1_address -> pio_key:address
	wire         mm_interconnect_0_pio_led_s1_chipselect;                     // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                       // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                        // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_write;                          // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                      // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire         mm_interconnect_0_sdram47_s1_chipselect;                     // mm_interconnect_0:sdram47_s1_chipselect -> sdram47:az_cs
	wire  [31:0] mm_interconnect_0_sdram47_s1_readdata;                       // sdram47:za_data -> mm_interconnect_0:sdram47_s1_readdata
	wire         mm_interconnect_0_sdram47_s1_waitrequest;                    // sdram47:za_waitrequest -> mm_interconnect_0:sdram47_s1_waitrequest
	wire  [20:0] mm_interconnect_0_sdram47_s1_address;                        // mm_interconnect_0:sdram47_s1_address -> sdram47:az_addr
	wire         mm_interconnect_0_sdram47_s1_read;                           // mm_interconnect_0:sdram47_s1_read -> sdram47:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram47_s1_byteenable;                     // mm_interconnect_0:sdram47_s1_byteenable -> sdram47:az_be_n
	wire         mm_interconnect_0_sdram47_s1_readdatavalid;                  // sdram47:za_valid -> mm_interconnect_0:sdram47_s1_readdatavalid
	wire         mm_interconnect_0_sdram47_s1_write;                          // mm_interconnect_0:sdram47_s1_write -> sdram47:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram47_s1_writedata;                      // mm_interconnect_0:sdram47_s1_writedata -> sdram47:az_data
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // epcs:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_irq_irq;                                               // irq_mapper:sender_irq -> nios2:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [epcs:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, pio_key:reset_n, pio_led:reset_n, ram:reset, rst_translator:in_reset, sdram47:reset_n, sysid_qsys_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [epcs:reset_req, nios2:reset_req, ram:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                             // nios2:debug_reset_request -> rst_controller:reset_in1

	nios2_qsys_epcs epcs (
		.clk        (clk_clk),                                             //               clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //             reset.reset_n
		.reset_req  (rst_controller_reset_out_reset_req),                  //                  .reset_req
		.address    (mm_interconnect_0_epcs_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_epcs_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_epcs_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_epcs_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_epcs_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_epcs_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_mapper_receiver1_irq),                            //               irq.irq
		.dclk       (epcs_dclk),                                           //          external.export
		.sce        (epcs_sce),                                            //                  .export
		.sdo        (epcs_sdo),                                            //                  .export
		.data0      (epcs_data0)                                           //                  .export
	);

	nios2_qsys_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios2_qsys_nios2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	nios2_qsys_pio_key pio_key (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_pio_key_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_key_s1_readdata), //                    .readdata
		.in_port  (key_export)                             // external_connection.export
	);

	nios2_qsys_pio_led pio_led (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                               // external_connection.export
	);

	nios2_qsys_ram ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	nios2_qsys_sdram47 sdram47 (
		.clk            (clk_clk),                                    //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),            // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram47_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram47_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram47_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram47_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram47_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram47_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram47_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram47_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram47_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram47_addr),                               //  wire.export
		.zs_ba          (sdram47_ba),                                 //      .export
		.zs_cas_n       (sdram47_cas_n),                              //      .export
		.zs_cke         (sdram47_cke),                                //      .export
		.zs_cs_n        (sdram47_cs_n),                               //      .export
		.zs_dq          (sdram47_dq),                                 //      .export
		.zs_dqm         (sdram47_dqm),                                //      .export
		.zs_ras_n       (sdram47_ras_n),                              //      .export
		.zs_we_n        (sdram47_we_n)                                //      .export
	);

	nios2_qsys_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios2_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                             (clk_clk),                                                     //                         clk_0_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                              // nios2_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address                 (nios2_data_master_address),                                   //                 nios2_data_master.address
		.nios2_data_master_waitrequest             (nios2_data_master_waitrequest),                               //                                  .waitrequest
		.nios2_data_master_byteenable              (nios2_data_master_byteenable),                                //                                  .byteenable
		.nios2_data_master_read                    (nios2_data_master_read),                                      //                                  .read
		.nios2_data_master_readdata                (nios2_data_master_readdata),                                  //                                  .readdata
		.nios2_data_master_readdatavalid           (nios2_data_master_readdatavalid),                             //                                  .readdatavalid
		.nios2_data_master_write                   (nios2_data_master_write),                                     //                                  .write
		.nios2_data_master_writedata               (nios2_data_master_writedata),                                 //                                  .writedata
		.nios2_data_master_debugaccess             (nios2_data_master_debugaccess),                               //                                  .debugaccess
		.nios2_instruction_master_address          (nios2_instruction_master_address),                            //          nios2_instruction_master.address
		.nios2_instruction_master_waitrequest      (nios2_instruction_master_waitrequest),                        //                                  .waitrequest
		.nios2_instruction_master_read             (nios2_instruction_master_read),                               //                                  .read
		.nios2_instruction_master_readdata         (nios2_instruction_master_readdata),                           //                                  .readdata
		.nios2_instruction_master_readdatavalid    (nios2_instruction_master_readdatavalid),                      //                                  .readdatavalid
		.epcs_epcs_control_port_address            (mm_interconnect_0_epcs_epcs_control_port_address),            //            epcs_epcs_control_port.address
		.epcs_epcs_control_port_write              (mm_interconnect_0_epcs_epcs_control_port_write),              //                                  .write
		.epcs_epcs_control_port_read               (mm_interconnect_0_epcs_epcs_control_port_read),               //                                  .read
		.epcs_epcs_control_port_readdata           (mm_interconnect_0_epcs_epcs_control_port_readdata),           //                                  .readdata
		.epcs_epcs_control_port_writedata          (mm_interconnect_0_epcs_epcs_control_port_writedata),          //                                  .writedata
		.epcs_epcs_control_port_chipselect         (mm_interconnect_0_epcs_epcs_control_port_chipselect),         //                                  .chipselect
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //     jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.nios2_debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),             //             nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),               //                                  .write
		.nios2_debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),                //                                  .read
		.nios2_debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),            //                                  .readdata
		.nios2_debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),           //                                  .writedata
		.nios2_debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),          //                                  .byteenable
		.nios2_debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),         //                                  .waitrequest
		.nios2_debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),         //                                  .debugaccess
		.pio_key_s1_address                        (mm_interconnect_0_pio_key_s1_address),                        //                        pio_key_s1.address
		.pio_key_s1_readdata                       (mm_interconnect_0_pio_key_s1_readdata),                       //                                  .readdata
		.pio_led_s1_address                        (mm_interconnect_0_pio_led_s1_address),                        //                        pio_led_s1.address
		.pio_led_s1_write                          (mm_interconnect_0_pio_led_s1_write),                          //                                  .write
		.pio_led_s1_readdata                       (mm_interconnect_0_pio_led_s1_readdata),                       //                                  .readdata
		.pio_led_s1_writedata                      (mm_interconnect_0_pio_led_s1_writedata),                      //                                  .writedata
		.pio_led_s1_chipselect                     (mm_interconnect_0_pio_led_s1_chipselect),                     //                                  .chipselect
		.ram_s1_address                            (mm_interconnect_0_ram_s1_address),                            //                            ram_s1.address
		.ram_s1_write                              (mm_interconnect_0_ram_s1_write),                              //                                  .write
		.ram_s1_readdata                           (mm_interconnect_0_ram_s1_readdata),                           //                                  .readdata
		.ram_s1_writedata                          (mm_interconnect_0_ram_s1_writedata),                          //                                  .writedata
		.ram_s1_byteenable                         (mm_interconnect_0_ram_s1_byteenable),                         //                                  .byteenable
		.ram_s1_chipselect                         (mm_interconnect_0_ram_s1_chipselect),                         //                                  .chipselect
		.ram_s1_clken                              (mm_interconnect_0_ram_s1_clken),                              //                                  .clken
		.sdram47_s1_address                        (mm_interconnect_0_sdram47_s1_address),                        //                        sdram47_s1.address
		.sdram47_s1_write                          (mm_interconnect_0_sdram47_s1_write),                          //                                  .write
		.sdram47_s1_read                           (mm_interconnect_0_sdram47_s1_read),                           //                                  .read
		.sdram47_s1_readdata                       (mm_interconnect_0_sdram47_s1_readdata),                       //                                  .readdata
		.sdram47_s1_writedata                      (mm_interconnect_0_sdram47_s1_writedata),                      //                                  .writedata
		.sdram47_s1_byteenable                     (mm_interconnect_0_sdram47_s1_byteenable),                     //                                  .byteenable
		.sdram47_s1_readdatavalid                  (mm_interconnect_0_sdram47_s1_readdatavalid),                  //                                  .readdatavalid
		.sdram47_s1_waitrequest                    (mm_interconnect_0_sdram47_s1_waitrequest),                    //                                  .waitrequest
		.sdram47_s1_chipselect                     (mm_interconnect_0_sdram47_s1_chipselect),                     //                                  .chipselect
		.sysid_qsys_0_control_slave_address        (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //        sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata       (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)        //                                  .readdata
	);

	nios2_qsys_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
